VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_wrapper
  CLASS BLOCK ;
  FOREIGN top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1700.000 ;
  PIN ADC_OUT_OBS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1472.920 1800.000 1473.520 ;
    END
  END ADC_OUT_OBS[0]
  PIN ADC_OUT_OBS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1562.000 1800.000 1562.600 ;
    END
  END ADC_OUT_OBS[1]
  PIN ADC_OUT_OBS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1651.080 1800.000 1651.680 ;
    END
  END ADC_OUT_OBS[2]
  PIN BL0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END BL0
  PIN CSA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 47.640 1800.000 48.240 ;
    END
  END CSA[0]
  PIN CSA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 938.440 1800.000 939.040 ;
    END
  END CSA[10]
  PIN CSA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1027.520 1800.000 1028.120 ;
    END
  END CSA[11]
  PIN CSA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1116.600 1800.000 1117.200 ;
    END
  END CSA[12]
  PIN CSA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1205.680 1800.000 1206.280 ;
    END
  END CSA[13]
  PIN CSA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1294.760 1800.000 1295.360 ;
    END
  END CSA[14]
  PIN CSA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1383.840 1800.000 1384.440 ;
    END
  END CSA[15]
  PIN CSA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 136.720 1800.000 137.320 ;
    END
  END CSA[1]
  PIN CSA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 225.800 1800.000 226.400 ;
    END
  END CSA[2]
  PIN CSA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 314.880 1800.000 315.480 ;
    END
  END CSA[3]
  PIN CSA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 403.960 1800.000 404.560 ;
    END
  END CSA[4]
  PIN CSA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 493.040 1800.000 493.640 ;
    END
  END CSA[5]
  PIN CSA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 582.120 1800.000 582.720 ;
    END
  END CSA[6]
  PIN CSA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 671.200 1800.000 671.800 ;
    END
  END CSA[7]
  PIN CSA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 760.280 1800.000 760.880 ;
    END
  END CSA[8]
  PIN CSA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 849.360 1800.000 849.960 ;
    END
  END CSA[9]
  PIN REF_CSA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.450 1696.000 1640.730 1700.000 ;
    END
  END REF_CSA
  PIN SL0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.830 0.000 1734.110 4.000 ;
    END
  END SL0
  PIN V0_REF_ADC
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 1696.000 1323.330 1700.000 ;
    END
  END V0_REF_ADC
  PIN V1_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1696.000 900.130 1700.000 ;
    END
  END V1_BL
  PIN V1_REF_ADC
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.850 1696.000 1429.130 1700.000 ;
    END
  END V1_REF_ADC
  PIN V1_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 1696.000 476.930 1700.000 ;
    END
  END V1_SL
  PIN V1_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 1696.000 53.730 1700.000 ;
    END
  END V1_WL
  PIN V2_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 1696.000 1005.930 1700.000 ;
    END
  END V2_BL
  PIN V2_REF_ADC
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 1696.000 1534.930 1700.000 ;
    END
  END V2_REF_ADC
  PIN V2_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 1696.000 582.730 1700.000 ;
    END
  END V2_SL
  PIN V2_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 1696.000 159.530 1700.000 ;
    END
  END V2_WL
  PIN V3_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 1696.000 1111.730 1700.000 ;
    END
  END V3_BL
  PIN V3_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 1696.000 688.530 1700.000 ;
    END
  END V3_SL
  PIN V3_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 1696.000 265.330 1700.000 ;
    END
  END V3_WL
  PIN V4_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1696.000 1217.530 1700.000 ;
    END
  END V4_BL
  PIN V4_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 1696.000 794.330 1700.000 ;
    END
  END V4_SL
  PIN V4_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 1696.000 371.130 1700.000 ;
    END
  END V4_WL
  PIN VDD_PRE
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.250 1696.000 1746.530 1700.000 ;
    END
  END VDD_PRE
  PIN WL0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 0.000 1751.130 4.000 ;
    END
  END WL0
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END clk
  PIN enable_IM
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END enable_IM
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 1696.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 1802.060 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 1695.120 1802.060 1696.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1800.460 3.280 1802.060 1696.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -0.020 22.640 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 -0.020 176.240 200.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 1107.725 176.240 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 -0.020 329.840 200.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 1107.725 329.840 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 -0.020 483.440 200.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 1107.725 483.440 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 -0.020 637.040 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 -0.020 790.640 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 1545.180 790.640 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 -0.020 944.240 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 1545.180 944.240 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 -0.020 1097.840 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 1545.180 1097.840 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 -0.020 1251.440 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 1545.180 1251.440 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 -0.020 1405.040 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 1545.180 1405.040 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 -0.020 1558.640 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 1545.180 1558.640 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 -0.020 1712.240 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 1545.180 1712.240 1700.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 26.730 1805.360 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 179.910 1805.360 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 333.090 688.340 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 486.270 688.340 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 639.450 688.340 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 792.630 688.340 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 945.810 688.340 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1098.990 688.340 1100.590 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1252.170 688.340 1253.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1405.350 688.340 1406.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1558.530 1805.360 1560.130 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 1700.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 1805.360 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1698.420 1805.360 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1803.760 -0.020 1805.360 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 -0.020 25.940 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 -0.020 179.540 200.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 1107.725 179.540 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 -0.020 333.140 200.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 1107.725 333.140 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 -0.020 486.740 200.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 1107.725 486.740 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 -0.020 640.340 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 -0.020 793.940 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 1545.180 793.940 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 -0.020 947.540 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 1545.180 947.540 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 -0.020 1101.140 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 1545.180 1101.140 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.140 -0.020 1254.740 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.140 1545.180 1254.740 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1406.740 -0.020 1408.340 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1406.740 1545.180 1408.340 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.340 -0.020 1561.940 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.340 1545.180 1561.940 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.940 -0.020 1715.540 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.940 1545.180 1715.540 1700.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 30.030 1805.360 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 183.210 1805.360 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 336.390 688.340 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 489.570 688.340 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 642.750 688.340 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 795.930 688.340 797.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 949.110 688.340 950.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1102.290 688.340 1103.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1255.470 688.340 1257.070 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1408.650 688.340 1410.250 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1561.830 1805.360 1563.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 217.360 601.100 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 239.120 601.100 261.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 266.320 601.100 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 315.280 601.100 326.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 331.600 601.100 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 386.000 601.100 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 402.320 601.100 430.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 456.720 601.100 468.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 478.480 601.100 500.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 527.440 601.100 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 549.200 601.100 571.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 598.160 601.100 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 619.920 601.100 642.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 668.880 601.100 680.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 690.640 601.100 701.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 701.745 601.100 712.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 739.600 601.100 750.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 761.360 601.100 783.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 599.500 810.320 601.100 821.680 ;
    END
  END vssd1
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END wbs_we_i
  PIN wishbone_address_bus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wishbone_address_bus[0]
  PIN wishbone_address_bus[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END wishbone_address_bus[10]
  PIN wishbone_address_bus[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END wishbone_address_bus[11]
  PIN wishbone_address_bus[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END wishbone_address_bus[12]
  PIN wishbone_address_bus[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END wishbone_address_bus[13]
  PIN wishbone_address_bus[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END wishbone_address_bus[14]
  PIN wishbone_address_bus[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END wishbone_address_bus[15]
  PIN wishbone_address_bus[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END wishbone_address_bus[16]
  PIN wishbone_address_bus[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END wishbone_address_bus[17]
  PIN wishbone_address_bus[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 0.000 1019.270 4.000 ;
    END
  END wishbone_address_bus[18]
  PIN wishbone_address_bus[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 0.000 1070.330 4.000 ;
    END
  END wishbone_address_bus[19]
  PIN wishbone_address_bus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wishbone_address_bus[1]
  PIN wishbone_address_bus[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END wishbone_address_bus[20]
  PIN wishbone_address_bus[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END wishbone_address_bus[21]
  PIN wishbone_address_bus[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 0.000 1223.510 4.000 ;
    END
  END wishbone_address_bus[22]
  PIN wishbone_address_bus[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END wishbone_address_bus[23]
  PIN wishbone_address_bus[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END wishbone_address_bus[24]
  PIN wishbone_address_bus[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.410 0.000 1376.690 4.000 ;
    END
  END wishbone_address_bus[25]
  PIN wishbone_address_bus[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.470 0.000 1427.750 4.000 ;
    END
  END wishbone_address_bus[26]
  PIN wishbone_address_bus[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 0.000 1478.810 4.000 ;
    END
  END wishbone_address_bus[27]
  PIN wishbone_address_bus[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END wishbone_address_bus[28]
  PIN wishbone_address_bus[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 0.000 1580.930 4.000 ;
    END
  END wishbone_address_bus[29]
  PIN wishbone_address_bus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wishbone_address_bus[2]
  PIN wishbone_address_bus[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.710 0.000 1631.990 4.000 ;
    END
  END wishbone_address_bus[30]
  PIN wishbone_address_bus[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.770 0.000 1683.050 4.000 ;
    END
  END wishbone_address_bus[31]
  PIN wishbone_address_bus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wishbone_address_bus[3]
  PIN wishbone_address_bus[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wishbone_address_bus[4]
  PIN wishbone_address_bus[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END wishbone_address_bus[5]
  PIN wishbone_address_bus[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END wishbone_address_bus[6]
  PIN wishbone_address_bus[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wishbone_address_bus[7]
  PIN wishbone_address_bus[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END wishbone_address_bus[8]
  PIN wishbone_address_bus[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END wishbone_address_bus[9]
  PIN wishbone_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wishbone_data_in[0]
  PIN wishbone_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wishbone_data_in[10]
  PIN wishbone_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END wishbone_data_in[11]
  PIN wishbone_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wishbone_data_in[12]
  PIN wishbone_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 4.000 ;
    END
  END wishbone_data_in[13]
  PIN wishbone_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END wishbone_data_in[14]
  PIN wishbone_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END wishbone_data_in[15]
  PIN wishbone_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END wishbone_data_in[16]
  PIN wishbone_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END wishbone_data_in[17]
  PIN wishbone_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END wishbone_data_in[18]
  PIN wishbone_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END wishbone_data_in[19]
  PIN wishbone_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wishbone_data_in[1]
  PIN wishbone_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END wishbone_data_in[20]
  PIN wishbone_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 4.000 ;
    END
  END wishbone_data_in[21]
  PIN wishbone_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 0.000 1240.530 4.000 ;
    END
  END wishbone_data_in[22]
  PIN wishbone_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END wishbone_data_in[23]
  PIN wishbone_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END wishbone_data_in[24]
  PIN wishbone_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 0.000 1393.710 4.000 ;
    END
  END wishbone_data_in[25]
  PIN wishbone_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 0.000 1444.770 4.000 ;
    END
  END wishbone_data_in[26]
  PIN wishbone_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 0.000 1495.830 4.000 ;
    END
  END wishbone_data_in[27]
  PIN wishbone_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.610 0.000 1546.890 4.000 ;
    END
  END wishbone_data_in[28]
  PIN wishbone_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END wishbone_data_in[29]
  PIN wishbone_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wishbone_data_in[2]
  PIN wishbone_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END wishbone_data_in[30]
  PIN wishbone_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.790 0.000 1700.070 4.000 ;
    END
  END wishbone_data_in[31]
  PIN wishbone_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wishbone_data_in[3]
  PIN wishbone_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END wishbone_data_in[4]
  PIN wishbone_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wishbone_data_in[5]
  PIN wishbone_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wishbone_data_in[6]
  PIN wishbone_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wishbone_data_in[7]
  PIN wishbone_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wishbone_data_in[8]
  PIN wishbone_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END wishbone_data_in[9]
  PIN wishbone_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wishbone_data_out[0]
  PIN wishbone_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END wishbone_data_out[10]
  PIN wishbone_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END wishbone_data_out[11]
  PIN wishbone_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END wishbone_data_out[12]
  PIN wishbone_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END wishbone_data_out[13]
  PIN wishbone_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END wishbone_data_out[14]
  PIN wishbone_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END wishbone_data_out[15]
  PIN wishbone_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END wishbone_data_out[16]
  PIN wishbone_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 0.000 1002.250 4.000 ;
    END
  END wishbone_data_out[17]
  PIN wishbone_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END wishbone_data_out[18]
  PIN wishbone_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END wishbone_data_out[19]
  PIN wishbone_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wishbone_data_out[1]
  PIN wishbone_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 4.000 ;
    END
  END wishbone_data_out[20]
  PIN wishbone_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 0.000 1206.490 4.000 ;
    END
  END wishbone_data_out[21]
  PIN wishbone_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END wishbone_data_out[22]
  PIN wishbone_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 4.000 ;
    END
  END wishbone_data_out[23]
  PIN wishbone_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 0.000 1359.670 4.000 ;
    END
  END wishbone_data_out[24]
  PIN wishbone_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END wishbone_data_out[25]
  PIN wishbone_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.510 0.000 1461.790 4.000 ;
    END
  END wishbone_data_out[26]
  PIN wishbone_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 0.000 1512.850 4.000 ;
    END
  END wishbone_data_out[27]
  PIN wishbone_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END wishbone_data_out[28]
  PIN wishbone_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 0.000 1614.970 4.000 ;
    END
  END wishbone_data_out[29]
  PIN wishbone_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wishbone_data_out[2]
  PIN wishbone_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.750 0.000 1666.030 4.000 ;
    END
  END wishbone_data_out[30]
  PIN wishbone_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 0.000 1717.090 4.000 ;
    END
  END wishbone_data_out[31]
  PIN wishbone_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wishbone_data_out[3]
  PIN wishbone_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wishbone_data_out[4]
  PIN wishbone_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wishbone_data_out[5]
  PIN wishbone_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wishbone_data_out[6]
  PIN wishbone_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END wishbone_data_out[7]
  PIN wishbone_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END wishbone_data_out[8]
  PIN wishbone_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END wishbone_data_out[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1794.460 1689.205 ;
      LAYER met1 ;
        RECT 5.520 6.840 1794.460 1689.360 ;
      LAYER met2 ;
        RECT 21.070 1695.720 53.170 1696.330 ;
        RECT 54.010 1695.720 158.970 1696.330 ;
        RECT 159.810 1695.720 264.770 1696.330 ;
        RECT 265.610 1695.720 370.570 1696.330 ;
        RECT 371.410 1695.720 476.370 1696.330 ;
        RECT 477.210 1695.720 582.170 1696.330 ;
        RECT 583.010 1695.720 687.970 1696.330 ;
        RECT 688.810 1695.720 793.770 1696.330 ;
        RECT 794.610 1695.720 899.570 1696.330 ;
        RECT 900.410 1695.720 1005.370 1696.330 ;
        RECT 1006.210 1695.720 1111.170 1696.330 ;
        RECT 1112.010 1695.720 1216.970 1696.330 ;
        RECT 1217.810 1695.720 1322.770 1696.330 ;
        RECT 1323.610 1695.720 1428.570 1696.330 ;
        RECT 1429.410 1695.720 1534.370 1696.330 ;
        RECT 1535.210 1695.720 1640.170 1696.330 ;
        RECT 1641.010 1695.720 1745.970 1696.330 ;
        RECT 1746.810 1695.720 1792.990 1696.330 ;
        RECT 21.070 4.280 1792.990 1695.720 ;
        RECT 21.070 4.000 31.550 4.280 ;
        RECT 32.390 4.000 48.570 4.280 ;
        RECT 49.410 4.000 65.590 4.280 ;
        RECT 66.430 4.000 82.610 4.280 ;
        RECT 83.450 4.000 99.630 4.280 ;
        RECT 100.470 4.000 116.650 4.280 ;
        RECT 117.490 4.000 133.670 4.280 ;
        RECT 134.510 4.000 150.690 4.280 ;
        RECT 151.530 4.000 167.710 4.280 ;
        RECT 168.550 4.000 184.730 4.280 ;
        RECT 185.570 4.000 201.750 4.280 ;
        RECT 202.590 4.000 218.770 4.280 ;
        RECT 219.610 4.000 235.790 4.280 ;
        RECT 236.630 4.000 252.810 4.280 ;
        RECT 253.650 4.000 269.830 4.280 ;
        RECT 270.670 4.000 286.850 4.280 ;
        RECT 287.690 4.000 303.870 4.280 ;
        RECT 304.710 4.000 320.890 4.280 ;
        RECT 321.730 4.000 337.910 4.280 ;
        RECT 338.750 4.000 354.930 4.280 ;
        RECT 355.770 4.000 371.950 4.280 ;
        RECT 372.790 4.000 388.970 4.280 ;
        RECT 389.810 4.000 405.990 4.280 ;
        RECT 406.830 4.000 423.010 4.280 ;
        RECT 423.850 4.000 440.030 4.280 ;
        RECT 440.870 4.000 457.050 4.280 ;
        RECT 457.890 4.000 474.070 4.280 ;
        RECT 474.910 4.000 491.090 4.280 ;
        RECT 491.930 4.000 508.110 4.280 ;
        RECT 508.950 4.000 525.130 4.280 ;
        RECT 525.970 4.000 542.150 4.280 ;
        RECT 542.990 4.000 559.170 4.280 ;
        RECT 560.010 4.000 576.190 4.280 ;
        RECT 577.030 4.000 593.210 4.280 ;
        RECT 594.050 4.000 610.230 4.280 ;
        RECT 611.070 4.000 627.250 4.280 ;
        RECT 628.090 4.000 644.270 4.280 ;
        RECT 645.110 4.000 661.290 4.280 ;
        RECT 662.130 4.000 678.310 4.280 ;
        RECT 679.150 4.000 695.330 4.280 ;
        RECT 696.170 4.000 712.350 4.280 ;
        RECT 713.190 4.000 729.370 4.280 ;
        RECT 730.210 4.000 746.390 4.280 ;
        RECT 747.230 4.000 763.410 4.280 ;
        RECT 764.250 4.000 780.430 4.280 ;
        RECT 781.270 4.000 797.450 4.280 ;
        RECT 798.290 4.000 814.470 4.280 ;
        RECT 815.310 4.000 831.490 4.280 ;
        RECT 832.330 4.000 848.510 4.280 ;
        RECT 849.350 4.000 865.530 4.280 ;
        RECT 866.370 4.000 882.550 4.280 ;
        RECT 883.390 4.000 899.570 4.280 ;
        RECT 900.410 4.000 916.590 4.280 ;
        RECT 917.430 4.000 933.610 4.280 ;
        RECT 934.450 4.000 950.630 4.280 ;
        RECT 951.470 4.000 967.650 4.280 ;
        RECT 968.490 4.000 984.670 4.280 ;
        RECT 985.510 4.000 1001.690 4.280 ;
        RECT 1002.530 4.000 1018.710 4.280 ;
        RECT 1019.550 4.000 1035.730 4.280 ;
        RECT 1036.570 4.000 1052.750 4.280 ;
        RECT 1053.590 4.000 1069.770 4.280 ;
        RECT 1070.610 4.000 1086.790 4.280 ;
        RECT 1087.630 4.000 1103.810 4.280 ;
        RECT 1104.650 4.000 1120.830 4.280 ;
        RECT 1121.670 4.000 1137.850 4.280 ;
        RECT 1138.690 4.000 1154.870 4.280 ;
        RECT 1155.710 4.000 1171.890 4.280 ;
        RECT 1172.730 4.000 1188.910 4.280 ;
        RECT 1189.750 4.000 1205.930 4.280 ;
        RECT 1206.770 4.000 1222.950 4.280 ;
        RECT 1223.790 4.000 1239.970 4.280 ;
        RECT 1240.810 4.000 1256.990 4.280 ;
        RECT 1257.830 4.000 1274.010 4.280 ;
        RECT 1274.850 4.000 1291.030 4.280 ;
        RECT 1291.870 4.000 1308.050 4.280 ;
        RECT 1308.890 4.000 1325.070 4.280 ;
        RECT 1325.910 4.000 1342.090 4.280 ;
        RECT 1342.930 4.000 1359.110 4.280 ;
        RECT 1359.950 4.000 1376.130 4.280 ;
        RECT 1376.970 4.000 1393.150 4.280 ;
        RECT 1393.990 4.000 1410.170 4.280 ;
        RECT 1411.010 4.000 1427.190 4.280 ;
        RECT 1428.030 4.000 1444.210 4.280 ;
        RECT 1445.050 4.000 1461.230 4.280 ;
        RECT 1462.070 4.000 1478.250 4.280 ;
        RECT 1479.090 4.000 1495.270 4.280 ;
        RECT 1496.110 4.000 1512.290 4.280 ;
        RECT 1513.130 4.000 1529.310 4.280 ;
        RECT 1530.150 4.000 1546.330 4.280 ;
        RECT 1547.170 4.000 1563.350 4.280 ;
        RECT 1564.190 4.000 1580.370 4.280 ;
        RECT 1581.210 4.000 1597.390 4.280 ;
        RECT 1598.230 4.000 1614.410 4.280 ;
        RECT 1615.250 4.000 1631.430 4.280 ;
        RECT 1632.270 4.000 1648.450 4.280 ;
        RECT 1649.290 4.000 1665.470 4.280 ;
        RECT 1666.310 4.000 1682.490 4.280 ;
        RECT 1683.330 4.000 1699.510 4.280 ;
        RECT 1700.350 4.000 1716.530 4.280 ;
        RECT 1717.370 4.000 1733.550 4.280 ;
        RECT 1734.390 4.000 1750.570 4.280 ;
        RECT 1751.410 4.000 1767.590 4.280 ;
        RECT 1768.430 4.000 1792.990 4.280 ;
      LAYER met3 ;
        RECT 21.050 1652.080 1796.450 1689.285 ;
        RECT 21.050 1650.680 1795.600 1652.080 ;
        RECT 21.050 1563.000 1796.450 1650.680 ;
        RECT 21.050 1561.600 1795.600 1563.000 ;
        RECT 21.050 1473.920 1796.450 1561.600 ;
        RECT 21.050 1472.520 1795.600 1473.920 ;
        RECT 21.050 1384.840 1796.450 1472.520 ;
        RECT 21.050 1383.440 1795.600 1384.840 ;
        RECT 21.050 1295.760 1796.450 1383.440 ;
        RECT 21.050 1294.360 1795.600 1295.760 ;
        RECT 21.050 1206.680 1796.450 1294.360 ;
        RECT 21.050 1205.280 1795.600 1206.680 ;
        RECT 21.050 1117.600 1796.450 1205.280 ;
        RECT 21.050 1116.200 1795.600 1117.600 ;
        RECT 21.050 1028.520 1796.450 1116.200 ;
        RECT 21.050 1027.120 1795.600 1028.520 ;
        RECT 21.050 939.440 1796.450 1027.120 ;
        RECT 21.050 938.040 1795.600 939.440 ;
        RECT 21.050 850.360 1796.450 938.040 ;
        RECT 21.050 848.960 1795.600 850.360 ;
        RECT 21.050 761.280 1796.450 848.960 ;
        RECT 21.050 759.880 1795.600 761.280 ;
        RECT 21.050 672.200 1796.450 759.880 ;
        RECT 21.050 670.800 1795.600 672.200 ;
        RECT 21.050 583.120 1796.450 670.800 ;
        RECT 21.050 581.720 1795.600 583.120 ;
        RECT 21.050 494.040 1796.450 581.720 ;
        RECT 21.050 492.640 1795.600 494.040 ;
        RECT 21.050 404.960 1796.450 492.640 ;
        RECT 21.050 403.560 1795.600 404.960 ;
        RECT 21.050 315.880 1796.450 403.560 ;
        RECT 21.050 314.480 1795.600 315.880 ;
        RECT 21.050 226.800 1796.450 314.480 ;
        RECT 21.050 225.400 1795.600 226.800 ;
        RECT 21.050 137.720 1796.450 225.400 ;
        RECT 21.050 136.320 1795.600 137.720 ;
        RECT 21.050 48.640 1796.450 136.320 ;
        RECT 21.050 47.240 1795.600 48.640 ;
        RECT 21.050 10.715 1796.450 47.240 ;
      LAYER met4 ;
        RECT 3.540 8.640 21.040 1690.860 ;
        RECT 22.640 8.640 24.340 1690.860 ;
        RECT 25.940 1107.725 174.640 1690.860 ;
        RECT 176.240 1107.725 177.940 1690.860 ;
        RECT 179.540 1107.725 328.240 1690.860 ;
        RECT 329.840 1107.725 331.540 1690.860 ;
        RECT 333.140 1107.725 481.840 1690.860 ;
        RECT 483.440 1107.725 485.140 1690.860 ;
        RECT 486.740 1107.725 635.440 1690.860 ;
        RECT 25.940 821.680 635.440 1107.725 ;
        RECT 25.940 810.320 599.500 821.680 ;
        RECT 601.100 810.320 635.440 821.680 ;
        RECT 25.940 783.600 635.440 810.320 ;
        RECT 25.940 761.360 599.500 783.600 ;
        RECT 601.100 761.360 635.440 783.600 ;
        RECT 25.940 750.960 635.440 761.360 ;
        RECT 25.940 739.600 599.500 750.960 ;
        RECT 601.100 739.600 635.440 750.960 ;
        RECT 25.940 712.880 635.440 739.600 ;
        RECT 25.940 701.745 599.500 712.880 ;
        RECT 601.100 701.745 635.440 712.880 ;
        RECT 25.940 701.520 635.440 701.745 ;
        RECT 25.940 690.640 599.500 701.520 ;
        RECT 601.100 690.640 635.440 701.520 ;
        RECT 25.940 680.240 635.440 690.640 ;
        RECT 25.940 668.880 599.500 680.240 ;
        RECT 601.100 668.880 635.440 680.240 ;
        RECT 25.940 642.160 635.440 668.880 ;
        RECT 25.940 619.920 599.500 642.160 ;
        RECT 601.100 619.920 635.440 642.160 ;
        RECT 25.940 609.520 635.440 619.920 ;
        RECT 25.940 598.160 599.500 609.520 ;
        RECT 601.100 598.160 635.440 609.520 ;
        RECT 25.940 571.440 635.440 598.160 ;
        RECT 25.940 549.200 599.500 571.440 ;
        RECT 601.100 549.200 635.440 571.440 ;
        RECT 25.940 538.800 635.440 549.200 ;
        RECT 25.940 527.440 599.500 538.800 ;
        RECT 601.100 527.440 635.440 538.800 ;
        RECT 25.940 500.720 635.440 527.440 ;
        RECT 25.940 478.480 599.500 500.720 ;
        RECT 601.100 478.480 635.440 500.720 ;
        RECT 25.940 468.080 635.440 478.480 ;
        RECT 25.940 456.720 599.500 468.080 ;
        RECT 601.100 456.720 635.440 468.080 ;
        RECT 25.940 430.000 635.440 456.720 ;
        RECT 25.940 402.320 599.500 430.000 ;
        RECT 601.100 402.320 635.440 430.000 ;
        RECT 25.940 397.360 635.440 402.320 ;
        RECT 25.940 386.000 599.500 397.360 ;
        RECT 601.100 386.000 635.440 397.360 ;
        RECT 25.940 359.280 635.440 386.000 ;
        RECT 25.940 331.600 599.500 359.280 ;
        RECT 601.100 331.600 635.440 359.280 ;
        RECT 25.940 326.640 635.440 331.600 ;
        RECT 25.940 315.280 599.500 326.640 ;
        RECT 601.100 315.280 635.440 326.640 ;
        RECT 25.940 288.560 635.440 315.280 ;
        RECT 25.940 266.320 599.500 288.560 ;
        RECT 601.100 266.320 635.440 288.560 ;
        RECT 25.940 261.360 635.440 266.320 ;
        RECT 25.940 239.120 599.500 261.360 ;
        RECT 601.100 239.120 635.440 261.360 ;
        RECT 25.940 228.720 635.440 239.120 ;
        RECT 25.940 217.360 599.500 228.720 ;
        RECT 601.100 217.360 635.440 228.720 ;
        RECT 25.940 200.755 635.440 217.360 ;
        RECT 25.940 8.640 174.640 200.755 ;
        RECT 176.240 8.640 177.940 200.755 ;
        RECT 179.540 8.640 328.240 200.755 ;
        RECT 329.840 8.640 331.540 200.755 ;
        RECT 333.140 8.640 481.840 200.755 ;
        RECT 483.440 8.640 485.140 200.755 ;
        RECT 486.740 8.640 635.440 200.755 ;
        RECT 637.040 8.640 638.740 1690.860 ;
        RECT 640.340 1545.180 789.040 1690.860 ;
        RECT 790.640 1545.180 792.340 1690.860 ;
        RECT 793.940 1545.180 942.640 1690.860 ;
        RECT 944.240 1545.180 945.940 1690.860 ;
        RECT 947.540 1545.180 1096.240 1690.860 ;
        RECT 1097.840 1545.180 1099.540 1690.860 ;
        RECT 1101.140 1545.180 1249.840 1690.860 ;
        RECT 1251.440 1545.180 1253.140 1690.860 ;
        RECT 1254.740 1545.180 1403.440 1690.860 ;
        RECT 1405.040 1545.180 1406.740 1690.860 ;
        RECT 1408.340 1545.180 1557.040 1690.860 ;
        RECT 1558.640 1545.180 1560.340 1690.860 ;
        RECT 1561.940 1545.180 1710.640 1690.860 ;
        RECT 1712.240 1545.180 1713.940 1690.860 ;
        RECT 1715.540 1545.180 1796.960 1690.860 ;
        RECT 640.340 206.780 1796.960 1545.180 ;
        RECT 640.340 8.640 789.040 206.780 ;
        RECT 790.640 8.640 792.340 206.780 ;
        RECT 793.940 8.640 942.640 206.780 ;
        RECT 944.240 8.640 945.940 206.780 ;
        RECT 947.540 8.640 1096.240 206.780 ;
        RECT 1097.840 8.640 1099.540 206.780 ;
        RECT 1101.140 8.640 1249.840 206.780 ;
        RECT 1251.440 8.640 1253.140 206.780 ;
        RECT 1254.740 8.640 1403.440 206.780 ;
        RECT 1405.040 8.640 1406.740 206.780 ;
        RECT 1408.340 8.640 1557.040 206.780 ;
        RECT 1558.640 8.640 1560.340 206.780 ;
        RECT 1561.940 8.640 1710.640 206.780 ;
        RECT 1712.240 8.640 1713.940 206.780 ;
        RECT 1715.540 8.640 1796.960 206.780 ;
      LAYER met5 ;
        RECT 3.540 1563.430 1796.960 1690.860 ;
        RECT 3.540 1560.130 1796.960 1561.830 ;
        RECT 3.540 1410.250 1796.960 1558.530 ;
        RECT 688.340 1408.650 1796.960 1410.250 ;
        RECT 3.540 1406.950 1796.960 1408.650 ;
        RECT 688.340 1405.350 1796.960 1406.950 ;
        RECT 3.540 1257.070 1796.960 1405.350 ;
        RECT 688.340 1255.470 1796.960 1257.070 ;
        RECT 3.540 1253.770 1796.960 1255.470 ;
        RECT 688.340 1252.170 1796.960 1253.770 ;
        RECT 3.540 1103.890 1796.960 1252.170 ;
        RECT 688.340 1102.290 1796.960 1103.890 ;
        RECT 3.540 1100.590 1796.960 1102.290 ;
        RECT 688.340 1098.990 1796.960 1100.590 ;
        RECT 3.540 950.710 1796.960 1098.990 ;
        RECT 688.340 949.110 1796.960 950.710 ;
        RECT 3.540 947.410 1796.960 949.110 ;
        RECT 688.340 945.810 1796.960 947.410 ;
        RECT 3.540 797.530 1796.960 945.810 ;
        RECT 688.340 795.930 1796.960 797.530 ;
        RECT 3.540 794.230 1796.960 795.930 ;
        RECT 688.340 792.630 1796.960 794.230 ;
        RECT 3.540 644.350 1796.960 792.630 ;
        RECT 688.340 642.750 1796.960 644.350 ;
        RECT 3.540 641.050 1796.960 642.750 ;
        RECT 688.340 639.450 1796.960 641.050 ;
        RECT 3.540 491.170 1796.960 639.450 ;
        RECT 688.340 489.570 1796.960 491.170 ;
        RECT 3.540 487.870 1796.960 489.570 ;
        RECT 688.340 486.270 1796.960 487.870 ;
        RECT 3.540 337.990 1796.960 486.270 ;
        RECT 688.340 336.390 1796.960 337.990 ;
        RECT 3.540 334.690 1796.960 336.390 ;
        RECT 688.340 333.090 1796.960 334.690 ;
        RECT 3.540 184.810 1796.960 333.090 ;
        RECT 3.540 181.510 1796.960 183.210 ;
        RECT 3.540 31.630 1796.960 179.910 ;
        RECT 3.540 28.330 1796.960 30.030 ;
        RECT 3.540 8.640 1796.960 26.730 ;
  END
END top_wrapper
END LIBRARY

