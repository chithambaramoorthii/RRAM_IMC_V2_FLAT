VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_wrapper
  CLASS BLOCK ;
  FOREIGN top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1700.000 ;
  PIN ADC_OUT_OBS[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1472.920 1800.000 1473.520 ;
    END
  END ADC_OUT_OBS[0]
  PIN ADC_OUT_OBS[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1562.000 1800.000 1562.600 ;
    END
  END ADC_OUT_OBS[1]
  PIN ADC_OUT_OBS[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1651.080 1800.000 1651.680 ;
    END
  END ADC_OUT_OBS[2]
  PIN BL0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END BL0
  PIN CSA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 47.640 1800.000 48.240 ;
    END
  END CSA[0]
  PIN CSA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 938.440 1800.000 939.040 ;
    END
  END CSA[10]
  PIN CSA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1027.520 1800.000 1028.120 ;
    END
  END CSA[11]
  PIN CSA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1116.600 1800.000 1117.200 ;
    END
  END CSA[12]
  PIN CSA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1205.680 1800.000 1206.280 ;
    END
  END CSA[13]
  PIN CSA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1294.760 1800.000 1295.360 ;
    END
  END CSA[14]
  PIN CSA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1383.840 1800.000 1384.440 ;
    END
  END CSA[15]
  PIN CSA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 136.720 1800.000 137.320 ;
    END
  END CSA[1]
  PIN CSA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 225.800 1800.000 226.400 ;
    END
  END CSA[2]
  PIN CSA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 314.880 1800.000 315.480 ;
    END
  END CSA[3]
  PIN CSA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 403.960 1800.000 404.560 ;
    END
  END CSA[4]
  PIN CSA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 493.040 1800.000 493.640 ;
    END
  END CSA[5]
  PIN CSA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 582.120 1800.000 582.720 ;
    END
  END CSA[6]
  PIN CSA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 671.200 1800.000 671.800 ;
    END
  END CSA[7]
  PIN CSA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 760.280 1800.000 760.880 ;
    END
  END CSA[8]
  PIN CSA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 849.360 1800.000 849.960 ;
    END
  END CSA[9]
  PIN REF_CSA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.450 1696.000 1640.730 1700.000 ;
    END
  END REF_CSA
  PIN SL0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.830 0.000 1734.110 4.000 ;
    END
  END SL0
  PIN V0_REF_ADC
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 1696.000 1323.330 1700.000 ;
    END
  END V0_REF_ADC
  PIN V1_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1696.000 900.130 1700.000 ;
    END
  END V1_BL
  PIN V1_REF_ADC
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.850 1696.000 1429.130 1700.000 ;
    END
  END V1_REF_ADC
  PIN V1_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 1696.000 476.930 1700.000 ;
    END
  END V1_SL
  PIN V1_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 1696.000 53.730 1700.000 ;
    END
  END V1_WL
  PIN V2_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 1696.000 1005.930 1700.000 ;
    END
  END V2_BL
  PIN V2_REF_ADC
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 1696.000 1534.930 1700.000 ;
    END
  END V2_REF_ADC
  PIN V2_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 1696.000 582.730 1700.000 ;
    END
  END V2_SL
  PIN V2_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 1696.000 159.530 1700.000 ;
    END
  END V2_WL
  PIN V3_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 1696.000 1111.730 1700.000 ;
    END
  END V3_BL
  PIN V3_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 1696.000 688.530 1700.000 ;
    END
  END V3_SL
  PIN V3_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 1696.000 265.330 1700.000 ;
    END
  END V3_WL
  PIN V4_BL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1696.000 1217.530 1700.000 ;
    END
  END V4_BL
  PIN V4_SL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 1696.000 794.330 1700.000 ;
    END
  END V4_SL
  PIN V4_WL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 1696.000 371.130 1700.000 ;
    END
  END V4_WL
  PIN VDD_PRE
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.250 1696.000 1746.530 1700.000 ;
    END
  END VDD_PRE
  PIN WL0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 0.000 1751.130 4.000 ;
    END
  END WL0
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END clk
  PIN enable_IM
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END enable_IM
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 1696.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 1802.060 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 1695.120 1802.060 1696.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1800.460 3.280 1802.060 1696.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -0.020 22.640 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 -0.020 176.240 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 -0.020 329.840 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 -0.020 483.440 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 -0.020 637.040 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 -0.020 790.640 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 1545.180 790.640 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 -0.020 944.240 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 1545.180 944.240 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 -0.020 1097.840 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 1545.180 1097.840 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 -0.020 1251.440 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 1545.180 1251.440 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 -0.020 1405.040 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 1545.180 1405.040 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 -0.020 1558.640 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 1545.180 1558.640 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 -0.020 1712.240 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 1545.180 1712.240 1700.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 26.730 1805.360 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 179.910 1805.360 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 333.090 688.340 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 486.270 688.340 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 639.450 688.340 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 792.630 688.340 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 945.810 688.340 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1098.990 688.340 1100.590 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1252.170 688.340 1253.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1405.350 688.340 1406.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1558.530 1805.360 1560.130 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 1700.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 1805.360 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1698.420 1805.360 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1803.760 -0.020 1805.360 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 -0.020 25.940 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 -0.020 179.540 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 -0.020 333.140 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 -0.020 486.740 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 -0.020 640.340 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 -0.020 793.940 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 1545.180 793.940 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 -0.020 947.540 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 1545.180 947.540 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 -0.020 1101.140 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 1545.180 1101.140 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.140 -0.020 1254.740 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.140 1545.180 1254.740 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1406.740 -0.020 1408.340 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1406.740 1545.180 1408.340 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.340 -0.020 1561.940 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.340 1545.180 1561.940 1700.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.940 -0.020 1715.540 206.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.940 1545.180 1715.540 1700.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 30.030 1805.360 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 183.210 1805.360 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 336.390 688.340 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 489.570 688.340 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 642.750 688.340 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 795.930 688.340 797.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 949.110 688.340 950.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1102.290 688.340 1103.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1255.470 688.340 1257.070 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1408.650 688.340 1410.250 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1561.830 1805.360 1563.430 ;
    END
  END vssd1
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END wbs_we_i
  PIN wishbone_address_bus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wishbone_address_bus[0]
  PIN wishbone_address_bus[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END wishbone_address_bus[10]
  PIN wishbone_address_bus[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END wishbone_address_bus[11]
  PIN wishbone_address_bus[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END wishbone_address_bus[12]
  PIN wishbone_address_bus[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END wishbone_address_bus[13]
  PIN wishbone_address_bus[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END wishbone_address_bus[14]
  PIN wishbone_address_bus[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END wishbone_address_bus[15]
  PIN wishbone_address_bus[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END wishbone_address_bus[16]
  PIN wishbone_address_bus[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END wishbone_address_bus[17]
  PIN wishbone_address_bus[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 0.000 1019.270 4.000 ;
    END
  END wishbone_address_bus[18]
  PIN wishbone_address_bus[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 0.000 1070.330 4.000 ;
    END
  END wishbone_address_bus[19]
  PIN wishbone_address_bus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wishbone_address_bus[1]
  PIN wishbone_address_bus[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END wishbone_address_bus[20]
  PIN wishbone_address_bus[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END wishbone_address_bus[21]
  PIN wishbone_address_bus[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 0.000 1223.510 4.000 ;
    END
  END wishbone_address_bus[22]
  PIN wishbone_address_bus[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END wishbone_address_bus[23]
  PIN wishbone_address_bus[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END wishbone_address_bus[24]
  PIN wishbone_address_bus[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.410 0.000 1376.690 4.000 ;
    END
  END wishbone_address_bus[25]
  PIN wishbone_address_bus[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.470 0.000 1427.750 4.000 ;
    END
  END wishbone_address_bus[26]
  PIN wishbone_address_bus[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 0.000 1478.810 4.000 ;
    END
  END wishbone_address_bus[27]
  PIN wishbone_address_bus[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END wishbone_address_bus[28]
  PIN wishbone_address_bus[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 0.000 1580.930 4.000 ;
    END
  END wishbone_address_bus[29]
  PIN wishbone_address_bus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wishbone_address_bus[2]
  PIN wishbone_address_bus[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.710 0.000 1631.990 4.000 ;
    END
  END wishbone_address_bus[30]
  PIN wishbone_address_bus[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.770 0.000 1683.050 4.000 ;
    END
  END wishbone_address_bus[31]
  PIN wishbone_address_bus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wishbone_address_bus[3]
  PIN wishbone_address_bus[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wishbone_address_bus[4]
  PIN wishbone_address_bus[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END wishbone_address_bus[5]
  PIN wishbone_address_bus[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END wishbone_address_bus[6]
  PIN wishbone_address_bus[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wishbone_address_bus[7]
  PIN wishbone_address_bus[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END wishbone_address_bus[8]
  PIN wishbone_address_bus[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END wishbone_address_bus[9]
  PIN wishbone_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wishbone_data_in[0]
  PIN wishbone_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wishbone_data_in[10]
  PIN wishbone_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END wishbone_data_in[11]
  PIN wishbone_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wishbone_data_in[12]
  PIN wishbone_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 4.000 ;
    END
  END wishbone_data_in[13]
  PIN wishbone_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END wishbone_data_in[14]
  PIN wishbone_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END wishbone_data_in[15]
  PIN wishbone_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END wishbone_data_in[16]
  PIN wishbone_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END wishbone_data_in[17]
  PIN wishbone_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END wishbone_data_in[18]
  PIN wishbone_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END wishbone_data_in[19]
  PIN wishbone_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wishbone_data_in[1]
  PIN wishbone_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END wishbone_data_in[20]
  PIN wishbone_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 4.000 ;
    END
  END wishbone_data_in[21]
  PIN wishbone_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 0.000 1240.530 4.000 ;
    END
  END wishbone_data_in[22]
  PIN wishbone_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END wishbone_data_in[23]
  PIN wishbone_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END wishbone_data_in[24]
  PIN wishbone_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 0.000 1393.710 4.000 ;
    END
  END wishbone_data_in[25]
  PIN wishbone_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 0.000 1444.770 4.000 ;
    END
  END wishbone_data_in[26]
  PIN wishbone_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 0.000 1495.830 4.000 ;
    END
  END wishbone_data_in[27]
  PIN wishbone_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.610 0.000 1546.890 4.000 ;
    END
  END wishbone_data_in[28]
  PIN wishbone_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END wishbone_data_in[29]
  PIN wishbone_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wishbone_data_in[2]
  PIN wishbone_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END wishbone_data_in[30]
  PIN wishbone_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.790 0.000 1700.070 4.000 ;
    END
  END wishbone_data_in[31]
  PIN wishbone_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wishbone_data_in[3]
  PIN wishbone_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END wishbone_data_in[4]
  PIN wishbone_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wishbone_data_in[5]
  PIN wishbone_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wishbone_data_in[6]
  PIN wishbone_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wishbone_data_in[7]
  PIN wishbone_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wishbone_data_in[8]
  PIN wishbone_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END wishbone_data_in[9]
  PIN wishbone_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wishbone_data_out[0]
  PIN wishbone_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END wishbone_data_out[10]
  PIN wishbone_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END wishbone_data_out[11]
  PIN wishbone_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END wishbone_data_out[12]
  PIN wishbone_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END wishbone_data_out[13]
  PIN wishbone_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END wishbone_data_out[14]
  PIN wishbone_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END wishbone_data_out[15]
  PIN wishbone_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END wishbone_data_out[16]
  PIN wishbone_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 0.000 1002.250 4.000 ;
    END
  END wishbone_data_out[17]
  PIN wishbone_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END wishbone_data_out[18]
  PIN wishbone_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END wishbone_data_out[19]
  PIN wishbone_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wishbone_data_out[1]
  PIN wishbone_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 4.000 ;
    END
  END wishbone_data_out[20]
  PIN wishbone_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 0.000 1206.490 4.000 ;
    END
  END wishbone_data_out[21]
  PIN wishbone_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END wishbone_data_out[22]
  PIN wishbone_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 4.000 ;
    END
  END wishbone_data_out[23]
  PIN wishbone_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 0.000 1359.670 4.000 ;
    END
  END wishbone_data_out[24]
  PIN wishbone_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END wishbone_data_out[25]
  PIN wishbone_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.510 0.000 1461.790 4.000 ;
    END
  END wishbone_data_out[26]
  PIN wishbone_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 0.000 1512.850 4.000 ;
    END
  END wishbone_data_out[27]
  PIN wishbone_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END wishbone_data_out[28]
  PIN wishbone_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 0.000 1614.970 4.000 ;
    END
  END wishbone_data_out[29]
  PIN wishbone_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wishbone_data_out[2]
  PIN wishbone_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.750 0.000 1666.030 4.000 ;
    END
  END wishbone_data_out[30]
  PIN wishbone_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 0.000 1717.090 4.000 ;
    END
  END wishbone_data_out[31]
  PIN wishbone_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wishbone_data_out[3]
  PIN wishbone_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wishbone_data_out[4]
  PIN wishbone_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wishbone_data_out[5]
  PIN wishbone_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wishbone_data_out[6]
  PIN wishbone_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END wishbone_data_out[7]
  PIN wishbone_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END wishbone_data_out[8]
  PIN wishbone_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END wishbone_data_out[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1794.460 1689.205 ;
      LAYER met1 ;
        RECT 5.520 6.500 1799.910 1689.360 ;
      LAYER met2 ;
        RECT 21.070 1695.720 53.170 1696.330 ;
        RECT 54.010 1695.720 158.970 1696.330 ;
        RECT 159.810 1695.720 264.770 1696.330 ;
        RECT 265.610 1695.720 370.570 1696.330 ;
        RECT 371.410 1695.720 476.370 1696.330 ;
        RECT 477.210 1695.720 582.170 1696.330 ;
        RECT 583.010 1695.720 687.970 1696.330 ;
        RECT 688.810 1695.720 793.770 1696.330 ;
        RECT 794.610 1695.720 899.570 1696.330 ;
        RECT 900.410 1695.720 1005.370 1696.330 ;
        RECT 1006.210 1695.720 1111.170 1696.330 ;
        RECT 1112.010 1695.720 1216.970 1696.330 ;
        RECT 1217.810 1695.720 1322.770 1696.330 ;
        RECT 1323.610 1695.720 1428.570 1696.330 ;
        RECT 1429.410 1695.720 1534.370 1696.330 ;
        RECT 1535.210 1695.720 1640.170 1696.330 ;
        RECT 1641.010 1695.720 1745.970 1696.330 ;
        RECT 1746.810 1695.720 1799.880 1696.330 ;
        RECT 21.070 4.280 1799.880 1695.720 ;
        RECT 21.070 3.670 31.550 4.280 ;
        RECT 32.390 3.670 48.570 4.280 ;
        RECT 49.410 3.670 65.590 4.280 ;
        RECT 66.430 3.670 82.610 4.280 ;
        RECT 83.450 3.670 99.630 4.280 ;
        RECT 100.470 3.670 116.650 4.280 ;
        RECT 117.490 3.670 133.670 4.280 ;
        RECT 134.510 3.670 150.690 4.280 ;
        RECT 151.530 3.670 167.710 4.280 ;
        RECT 168.550 3.670 184.730 4.280 ;
        RECT 185.570 3.670 201.750 4.280 ;
        RECT 202.590 3.670 218.770 4.280 ;
        RECT 219.610 3.670 235.790 4.280 ;
        RECT 236.630 3.670 252.810 4.280 ;
        RECT 253.650 3.670 269.830 4.280 ;
        RECT 270.670 3.670 286.850 4.280 ;
        RECT 287.690 3.670 303.870 4.280 ;
        RECT 304.710 3.670 320.890 4.280 ;
        RECT 321.730 3.670 337.910 4.280 ;
        RECT 338.750 3.670 354.930 4.280 ;
        RECT 355.770 3.670 371.950 4.280 ;
        RECT 372.790 3.670 388.970 4.280 ;
        RECT 389.810 3.670 405.990 4.280 ;
        RECT 406.830 3.670 423.010 4.280 ;
        RECT 423.850 3.670 440.030 4.280 ;
        RECT 440.870 3.670 457.050 4.280 ;
        RECT 457.890 3.670 474.070 4.280 ;
        RECT 474.910 3.670 491.090 4.280 ;
        RECT 491.930 3.670 508.110 4.280 ;
        RECT 508.950 3.670 525.130 4.280 ;
        RECT 525.970 3.670 542.150 4.280 ;
        RECT 542.990 3.670 559.170 4.280 ;
        RECT 560.010 3.670 576.190 4.280 ;
        RECT 577.030 3.670 593.210 4.280 ;
        RECT 594.050 3.670 610.230 4.280 ;
        RECT 611.070 3.670 627.250 4.280 ;
        RECT 628.090 3.670 644.270 4.280 ;
        RECT 645.110 3.670 661.290 4.280 ;
        RECT 662.130 3.670 678.310 4.280 ;
        RECT 679.150 3.670 695.330 4.280 ;
        RECT 696.170 3.670 712.350 4.280 ;
        RECT 713.190 3.670 729.370 4.280 ;
        RECT 730.210 3.670 746.390 4.280 ;
        RECT 747.230 3.670 763.410 4.280 ;
        RECT 764.250 3.670 780.430 4.280 ;
        RECT 781.270 3.670 797.450 4.280 ;
        RECT 798.290 3.670 814.470 4.280 ;
        RECT 815.310 3.670 831.490 4.280 ;
        RECT 832.330 3.670 848.510 4.280 ;
        RECT 849.350 3.670 865.530 4.280 ;
        RECT 866.370 3.670 882.550 4.280 ;
        RECT 883.390 3.670 899.570 4.280 ;
        RECT 900.410 3.670 916.590 4.280 ;
        RECT 917.430 3.670 933.610 4.280 ;
        RECT 934.450 3.670 950.630 4.280 ;
        RECT 951.470 3.670 967.650 4.280 ;
        RECT 968.490 3.670 984.670 4.280 ;
        RECT 985.510 3.670 1001.690 4.280 ;
        RECT 1002.530 3.670 1018.710 4.280 ;
        RECT 1019.550 3.670 1035.730 4.280 ;
        RECT 1036.570 3.670 1052.750 4.280 ;
        RECT 1053.590 3.670 1069.770 4.280 ;
        RECT 1070.610 3.670 1086.790 4.280 ;
        RECT 1087.630 3.670 1103.810 4.280 ;
        RECT 1104.650 3.670 1120.830 4.280 ;
        RECT 1121.670 3.670 1137.850 4.280 ;
        RECT 1138.690 3.670 1154.870 4.280 ;
        RECT 1155.710 3.670 1171.890 4.280 ;
        RECT 1172.730 3.670 1188.910 4.280 ;
        RECT 1189.750 3.670 1205.930 4.280 ;
        RECT 1206.770 3.670 1222.950 4.280 ;
        RECT 1223.790 3.670 1239.970 4.280 ;
        RECT 1240.810 3.670 1256.990 4.280 ;
        RECT 1257.830 3.670 1274.010 4.280 ;
        RECT 1274.850 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1308.050 4.280 ;
        RECT 1308.890 3.670 1325.070 4.280 ;
        RECT 1325.910 3.670 1342.090 4.280 ;
        RECT 1342.930 3.670 1359.110 4.280 ;
        RECT 1359.950 3.670 1376.130 4.280 ;
        RECT 1376.970 3.670 1393.150 4.280 ;
        RECT 1393.990 3.670 1410.170 4.280 ;
        RECT 1411.010 3.670 1427.190 4.280 ;
        RECT 1428.030 3.670 1444.210 4.280 ;
        RECT 1445.050 3.670 1461.230 4.280 ;
        RECT 1462.070 3.670 1478.250 4.280 ;
        RECT 1479.090 3.670 1495.270 4.280 ;
        RECT 1496.110 3.670 1512.290 4.280 ;
        RECT 1513.130 3.670 1529.310 4.280 ;
        RECT 1530.150 3.670 1546.330 4.280 ;
        RECT 1547.170 3.670 1563.350 4.280 ;
        RECT 1564.190 3.670 1580.370 4.280 ;
        RECT 1581.210 3.670 1597.390 4.280 ;
        RECT 1598.230 3.670 1614.410 4.280 ;
        RECT 1615.250 3.670 1631.430 4.280 ;
        RECT 1632.270 3.670 1648.450 4.280 ;
        RECT 1649.290 3.670 1665.470 4.280 ;
        RECT 1666.310 3.670 1682.490 4.280 ;
        RECT 1683.330 3.670 1699.510 4.280 ;
        RECT 1700.350 3.670 1716.530 4.280 ;
        RECT 1717.370 3.670 1733.550 4.280 ;
        RECT 1734.390 3.670 1750.570 4.280 ;
        RECT 1751.410 3.670 1767.590 4.280 ;
        RECT 1768.430 3.670 1799.880 4.280 ;
      LAYER met3 ;
        RECT 21.050 1652.080 1796.235 1689.285 ;
        RECT 21.050 1650.680 1795.600 1652.080 ;
        RECT 21.050 1563.000 1796.235 1650.680 ;
        RECT 21.050 1561.600 1795.600 1563.000 ;
        RECT 21.050 1473.920 1796.235 1561.600 ;
        RECT 21.050 1472.520 1795.600 1473.920 ;
        RECT 21.050 1384.840 1796.235 1472.520 ;
        RECT 21.050 1383.440 1795.600 1384.840 ;
        RECT 21.050 1295.760 1796.235 1383.440 ;
        RECT 21.050 1294.360 1795.600 1295.760 ;
        RECT 21.050 1206.680 1796.235 1294.360 ;
        RECT 21.050 1205.280 1795.600 1206.680 ;
        RECT 21.050 1117.600 1796.235 1205.280 ;
        RECT 21.050 1116.200 1795.600 1117.600 ;
        RECT 21.050 1028.520 1796.235 1116.200 ;
        RECT 21.050 1027.120 1795.600 1028.520 ;
        RECT 21.050 939.440 1796.235 1027.120 ;
        RECT 21.050 938.040 1795.600 939.440 ;
        RECT 21.050 850.360 1796.235 938.040 ;
        RECT 21.050 848.960 1795.600 850.360 ;
        RECT 21.050 761.280 1796.235 848.960 ;
        RECT 21.050 759.880 1795.600 761.280 ;
        RECT 21.050 672.200 1796.235 759.880 ;
        RECT 21.050 670.800 1795.600 672.200 ;
        RECT 21.050 583.120 1796.235 670.800 ;
        RECT 21.050 581.720 1795.600 583.120 ;
        RECT 21.050 494.040 1796.235 581.720 ;
        RECT 21.050 492.640 1795.600 494.040 ;
        RECT 21.050 404.960 1796.235 492.640 ;
        RECT 21.050 403.560 1795.600 404.960 ;
        RECT 21.050 315.880 1796.235 403.560 ;
        RECT 21.050 314.480 1795.600 315.880 ;
        RECT 21.050 226.800 1796.235 314.480 ;
        RECT 21.050 225.400 1795.600 226.800 ;
        RECT 21.050 137.720 1796.235 225.400 ;
        RECT 21.050 136.320 1795.600 137.720 ;
        RECT 21.050 48.640 1796.235 136.320 ;
        RECT 21.050 47.240 1795.600 48.640 ;
        RECT 21.050 8.335 1796.235 47.240 ;
      LAYER met4 ;
        RECT 242.255 11.735 327.840 1622.305 ;
        RECT 330.240 11.735 331.140 1622.305 ;
        RECT 333.540 11.735 481.440 1622.305 ;
        RECT 483.840 11.735 484.740 1622.305 ;
        RECT 487.140 11.735 635.040 1622.305 ;
        RECT 637.440 11.735 638.340 1622.305 ;
        RECT 640.740 1544.780 788.640 1622.305 ;
        RECT 791.040 1544.780 791.940 1622.305 ;
        RECT 794.340 1544.780 942.240 1622.305 ;
        RECT 944.640 1544.780 945.540 1622.305 ;
        RECT 947.940 1544.780 1095.840 1622.305 ;
        RECT 1098.240 1544.780 1099.140 1622.305 ;
        RECT 1101.540 1544.780 1249.440 1622.305 ;
        RECT 1251.840 1544.780 1252.740 1622.305 ;
        RECT 1255.140 1544.780 1403.040 1622.305 ;
        RECT 1405.440 1544.780 1406.340 1622.305 ;
        RECT 1408.740 1544.780 1556.640 1622.305 ;
        RECT 1559.040 1544.780 1559.940 1622.305 ;
        RECT 1562.340 1544.780 1710.240 1622.305 ;
        RECT 1712.640 1544.780 1713.540 1622.305 ;
        RECT 1715.940 1544.780 1789.105 1622.305 ;
        RECT 640.740 207.180 1789.105 1544.780 ;
        RECT 640.740 11.735 788.640 207.180 ;
        RECT 791.040 11.735 791.940 207.180 ;
        RECT 794.340 11.735 942.240 207.180 ;
        RECT 944.640 11.735 945.540 207.180 ;
        RECT 947.940 11.735 1095.840 207.180 ;
        RECT 1098.240 11.735 1099.140 207.180 ;
        RECT 1101.540 11.735 1249.440 207.180 ;
        RECT 1251.840 11.735 1252.740 207.180 ;
        RECT 1255.140 11.735 1403.040 207.180 ;
        RECT 1405.440 11.735 1406.340 207.180 ;
        RECT 1408.740 11.735 1556.640 207.180 ;
        RECT 1559.040 11.735 1559.940 207.180 ;
        RECT 1562.340 11.735 1710.240 207.180 ;
        RECT 1712.640 11.735 1713.540 207.180 ;
        RECT 1715.940 11.735 1789.105 207.180 ;
      LAYER met5 ;
        RECT 657.770 1411.850 1756.280 1534.880 ;
        RECT 689.940 1403.750 1756.280 1411.850 ;
        RECT 657.770 1258.670 1756.280 1403.750 ;
        RECT 689.940 1250.570 1756.280 1258.670 ;
        RECT 657.770 1105.490 1756.280 1250.570 ;
        RECT 689.940 1097.390 1756.280 1105.490 ;
        RECT 657.770 952.310 1756.280 1097.390 ;
        RECT 689.940 944.210 1756.280 952.310 ;
        RECT 657.770 799.130 1756.280 944.210 ;
        RECT 689.940 791.030 1756.280 799.130 ;
        RECT 657.770 645.950 1756.280 791.030 ;
        RECT 689.940 637.850 1756.280 645.950 ;
        RECT 657.770 492.770 1756.280 637.850 ;
        RECT 689.940 484.670 1756.280 492.770 ;
        RECT 657.770 339.590 1756.280 484.670 ;
        RECT 689.940 331.490 1756.280 339.590 ;
        RECT 657.770 217.080 1756.280 331.490 ;
  END
END top_wrapper
END LIBRARY

